module data_ram(
    input wire clk,
    input wire rst,
    
    input wire we_i,
    input wire[31:0] addr_i,
    input wire[31:0] data_i,
    
    output reg[31:0] data_o
);
    
    reg[31:0] _ram[0:120071];
    integer i;
    initial begin
		_ram[16747] = 32'h00626261;
		_ram[16748] = 32'h00756f79;
		_ram[16749] = 32'h00746f6e;
		_ram[16750] = 32'h00007469;
		_ram[16751] = 32'h00646164;
		_ram[16752] = 32'h62626163;
		_ram[16753] = 32'h00006569;
		_ram[16754] = 32'h72756f79;
		_ram[16755] = 32'h00000000;
		_ram[16756] = 32'h69207449;
		_ram[16757] = 32'h74276e73;
		_ram[16758] = 32'h72656820;
		_ram[16759] = 32'h00000065;
		_ram[16760] = 32'h20747542;
		_ram[16761] = 32'h69207469;
		_ram[16762] = 32'h65682073;
		_ram[16763] = 32'h00006572;
		_ram[16764] = 32'h61646f68;
		_ram[16765] = 32'h00000064;
		_ram[16766] = 32'h686f6f79;
		_ram[16767] = 32'h00006f6f;
		_ram[16768] = 32'h00007878;
		_ram[16769] = 32'h00000078;
		_ram[16770] = 32'h0000002e;
		_ram[16771] = 32'h72206e49;
		_ram[16772] = 32'h6e656365;
		_ram[16773] = 32'h65792074;
		_ram[16774] = 32'h2c737261;
		_ram[16775] = 32'h65687420;
		_ram[16776] = 32'h65696620;
		_ram[16777] = 32'h6f20646c;
		_ram[16778] = 32'h68702066;
		_ram[16779] = 32'h6e6f746f;
		_ram[16780] = 32'h00206369;
		_ram[16781] = 32'h73797263;
		_ram[16782] = 32'h736c6174;
		_ram[16783] = 32'h73616820;
		_ram[16784] = 32'h756f6620;
		_ram[16785] = 32'h6e20646e;
		_ram[16786] = 32'h00007765;
		_ram[16787] = 32'h000105ac;
		_ram[16788] = 32'h000105b0;
		_ram[16789] = 32'h000105b4;
		_ram[16790] = 32'h000105b8;
		_ram[16791] = 32'h000105bc;
		_ram[16792] = 32'h00000000;
		_ram[16793] = 32'h000105c0;
		_ram[16794] = 32'h000105c8;
		_ram[16795] = 32'h000105d0;
		_ram[16796] = 32'h000105e0;
		_ram[16797] = 32'h000105f0;
		_ram[16798] = 32'h000105f8;
		_ram[16799] = 32'h000105f8;
		_ram[16800] = 32'h000105f8;
		_ram[16801] = 32'h000105f8;
		_ram[16802] = 32'h000105f8;
		_ram[16803] = 32'h00010600;
		_ram[16804] = 32'h00010604;
		_ram[16805] = 32'h00010608;
		_ram[16806] = 32'h0001060c;
		_ram[16807] = 32'h00010634;
		for(i=18436;i<18700;i=i+1)begin
		  _ram[i] = 0;
		end
		_ram[16357] = 32'h000105c0;
		_ram[16358] = 32'h000105c8;
    end
    always @ (posedge clk)begin
        if(we_i)begin
            _ram[addr_i[31:2]] <= data_i;
            
        end
    end
    
    always @ (*)begin
        if(rst)begin
            data_o = 0;
        end else begin
            data_o = _ram[addr_i[31:2]];
        end
    end
endmodule